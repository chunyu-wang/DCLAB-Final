module RGB2GRAY(
    input i_clk,
    input i_rst_n,
    input 
)



endmodule