`timescale 1ps/1ps

module testBackgroundSub(

);
    BackgroundSub(

    );
endmodule